{
"130":[0.5,1,0,2,8,8,300,0],
"131":[0.5,1,0,2,8,8,300,0],
"132":[0.5,1,0,2,8,8,300,0],
"133":[0.5,1,0,2,8,8,300,0],
"134":[0.5,1,0,2,8,8,300,0]
}