{
"ATTACK_COOLDOWN": 0.5,
"ATTACK_DMG": 1,
"ATTACK_EFFECT": 0,
"ATTACK_STACK": 2,
"CHAR_CODE": 130,
"HP": 10,
"MAX_HP": 10,
"MAX_SPEED": 300,
"SPECIAL_CODE": 0
}